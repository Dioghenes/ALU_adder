library ieee;
use ieee.std_logic_1164.all;

entity P4ADD is
		generic(log2_N_BIT: integer := 5);
		port(	A	    : in std_logic_vector(2**log2_N_BIT-1 downto 0);
			 	B 	    : in std_logic_vector(2**log2_N_BIT-1 downto 0);
				AddSub  : in std_logic;
				SUM     : out std_logic_vector(2**log2_N_BIT-1 downto 0);
			 	Cout	: out std_logic);
end entity;

architecture structural of P4ADD is
	
	-- Used component
	component sparsetree_radix4 is
		generic(log2_N_BIT : integer := 5);
		port(A	 : in std_logic_vector(2**log2_N_BIT-1 downto 0);		-- Operand A
			 B   : in std_logic_vector(2**log2_N_BIT-1 downto 0);		-- Operand B
			 Cin : in std_logic;										-- First carry in
			 g_o : out std_logic_vector((2**log2_N_BIT)/4 downto 0));	-- Carry vector generated
	end component;
	
	component sum_generator is
		generic(log2_N_BIT : integer := 5);
		port(A	  : in std_logic_vector(2**log2_N_BIT-1 downto 0);
			 B     : in std_logic_vector(2**log2_N_BIT-1 downto 0);
			 Cin   : in std_logic_vector((2**log2_N_BIT)/4-1 downto 0);
			 SUM   : out std_logic_vector(2**log2_N_BIT-1 downto 0));
	end component;
	
	-- Internal signals
	signal gout_sig : std_logic_vector((2**log2_N_BIT)/4 downto 0);
	signal B_int    : std_logic_vector(2**log2_N_BIT-1 downto 0);
	
begin
	-- XOR wall used to perform ADD or SUB according to AddSub signal
	XOR_gen : for i in 0 to 2**log2_N_BIT-1 generate
		B_int(i) <= B(i) xor AddSub; 
	end generate XOR_gen;
	
	-- Sparse tree carry generator
	ST : sparsetree_radix4 generic map(log2_N_BIT)
						   port map(A, B_int, AddSub, gout_sig);
								  
	-- Sum generator
	SG : sum_generator 	generic map(log2_N_BIT)
					    port map(A, B_int, gout_sig((2**log2_N_BIT)/4-1 downto 0), SUM);
	
	-- Cout generated by the sparse tree 
	Cout <= gout_sig((2**log2_N_BIT)/4);
	
end architecture;
